[aimspice]
[description]
629
CMOS_TSL
.subckt NOT_CMOS i vdd vss out
mn out i vss vss nmos1 l=1u w=1u
.model nmos1 nmos vto=1.5
mp out i vdd vdd pmos1 l=1u w=1u
.model pmos1 pmos vto=-1.5
.ends

.subckt NOT_CMOS_TSL in e vdd vss out
mn 2 e vss vss nmos1 l=1u w=1u
.model nmos1 nmos vto=1.5
mp 1 note vdd vdd pmos1 l=1u w=1u
.model pmos1 pmos vto=-1.5
X1_NOT_CMOS in 1 2 out NOT_CMOS
X2_NOT_CMOS e vdd vss note NOT_CMOS
.ends
X3_NOT_CMOS_TSL in e vdd vss out NOT_CMOS_TSL
R1 vdd out 1e6
R2 out vss 1e6
Cs1 out 0 15p
vdd vdd 0 5
vss vss 0 0
vi in 0 dc 5 pulse(0.1 4.8 0 1e-9 1e-9 1e-3 2e-3)
ve e 0 dc 0 pulse(0.2 4.9 1e-9 1e-9 2e-3 4e-3)
[dc]
1
vi
-1
5
0.01
[tran]
1e-2
5e-3
X
X
0
[ana]
1 1
0
1 1
1 1 -2 6
3
v(e)
v(out)
v(in)
[end]
