[aimspice]
[description]
210
redresor cu filtru
.Model Dioda D
D1 1 2 Dioda
D2 0 1 Dioda
D3 0 3 Dioda
D4 3 2 Dioda
R1 2 0 100
c1 2 0 30m
Vin 1 3 sin(0 10 1k 0 0)

!aduce din c.a. in c.c astfel si pe grafic obtinem o linie dreapta
[tran]
1e-9
6e-3
0
0.0001
0
[ana]
4 5
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
0
1 1
1 1 0 5
3
v(1)
v(2)
v(3)
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
0
1 1
1 1 -2 10
2
v(1)
v(2)
0
1 1
1 1 -2 10
2
v(1)
v(2)
[end]
