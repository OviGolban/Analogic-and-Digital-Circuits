[aimspice]
[description]
134
redresor dublaalternanta
.Model Dioda D
D1 1 2 Dioda
D2 0 1 Dioda
D3 0 3 Dioda
D4 3 2 Dioda
R1 2 0 100
Vin 1 3 sin(0 10 1k 0 0)
[tran]
1e-9
6e-3
0
0.0001
0
[ana]
4 1
0
1 1
1 1 -2 10
2
v(1)
v(2)
[end]
