[aimspice]
[description]
348
stabilizator parametric cu dioda zener
.Model Dioda D
.model zener d bv = 5.6
D1 1 2 Dioda
D2 0 1 Dioda
D3 0 3 Dioda
D4 3 2 Dioda
R1 2 0 100
c1 2 0 1m
dz 0 2 zener
Vin 1 3 sin(0 10 1k 0 0)

!dioda consuma o parte din curent, astfel observam ca  amplitudinea tensiunii este mai mcia decat in cazul in care am scoate dioda din circuit


[tran]
1e-9
6e-3
0
0.0001
0
[ana]
4 9
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
0
1 1
1 1 -80 20
4
v(1)
v(2)
v(3)
i(vin)
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
0
1 1
1 1 -2 10
2
v(1)
v(2)
0
1 1
1 1 -2 10
2
v(1)
v(2)
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
0
1 1
1 1 0 5
3
v(1)
v(2)
v(3)
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
[end]
